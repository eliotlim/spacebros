../../clarvi_fpga/prescale_int.sv