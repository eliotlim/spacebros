../../clarvi_fpga/prescale_pwr.sv